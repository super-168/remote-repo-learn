//  Class: Untitled-1
//
class Untitled-1;
    //  Group: Variables


    //  Group: Constraints


    //  Group: Functions

    //  Constructor: new
    function new(string name = "Untitled-1");
    endfunction: new
    

endclass: Untitled-1
