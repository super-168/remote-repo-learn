always_comb begin: <process_label>
    
end: <process_label>